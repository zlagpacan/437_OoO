`ifndef PRINT_MACROS_VH
`define PRINT_MACROS_VH

`define INFO_PRINTS
`define ERROR_PRINTS

`endif